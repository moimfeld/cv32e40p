VFADD_S            = 32'b1000001??????????000?????0110011
VFADD_R_S          = 32'b1000001??????????100?????0110011
VFSUB_S            = 32'b1000010??????????000?????0110011
VFSUB_R_S          = 32'b1000010??????????100?????0110011
VFMUL_S            = 32'b1000011??????????000?????0110011
VFMUL_R_S          = 32'b1000011??????????100?????0110011
VFDIV_S            = 32'b1000100??????????000?????0110011
VFDIV_R_S          = 32'b1000100??????????100?????0110011
VFMIN_S            = 32'b1000101??????????000?????0110011
VFMIN_R_S          = 32'b1000101??????????100?????0110011
VFMAX_S            = 32'b1000110??????????000?????0110011
VFMAX_R_S          = 32'b1000110??????????100?????0110011
VFSQRT_S           = 32'b100011100000?????000?????0110011
VFMAC_S            = 32'b1001000??????????000?????0110011
VFMAC_R_S          = 32'b1001000??????????100?????0110011
VFMRE_S            = 32'b1001001??????????000?????0110011
VFMRE_R_S          = 32'b1001001??????????100?????0110011
VFCLASS_S          = 32'b100110000001?????000?????0110011
VFSGNJ_S           = 32'b1001101??????????000?????0110011
VFSGNJ_R_S         = 32'b1001101??????????100?????0110011
VFSGNJN_S          = 32'b1001110??????????000?????0110011
VFSGNJN_R_S        = 32'b1001110??????????100?????0110011
VFSGNJX_S          = 32'b1001111??????????000?????0110011
VFSGNJX_R_S        = 32'b1001111??????????100?????0110011
VFEQ_S             = 32'b1010000??????????000?????0110011
VFEQ_R_S           = 32'b1010000??????????100?????0110011
VFNE_S             = 32'b1010001??????????000?????0110011
VFNE_R_S           = 32'b1010001??????????100?????0110011
VFLT_S             = 32'b1010010??????????000?????0110011
VFLT_R_S           = 32'b1010010??????????100?????0110011
VFGE_S             = 32'b1010011??????????000?????0110011
VFGE_R_S           = 32'b1010011??????????100?????0110011
VFLE_S             = 32'b1010100??????????000?????0110011
VFLE_R_S           = 32'b1010100??????????100?????0110011
VFGT_S             = 32'b1010101??????????000?????0110011
VFGT_R_S           = 32'b1010101??????????100?????0110011
VFMV_X_S           = 32'b100110000000?????000?????0110011
VFMV_S_X           = 32'b100110000000?????100?????0110011
VFCVT_X_S          = 32'b100110000010?????000?????0110011
VFCVT_XU_S         = 32'b100110000010?????100?????0110011
VFCVT_S_X          = 32'b100110000011?????000?????0110011
VFCVT_S_XU         = 32'b100110000011?????100?????0110011
VFCPKA_S_S         = 32'b1011000??????????000?????0110011
VFCPKB_S_S         = 32'b1011000??????????100?????0110011
VFCPKC_S_S         = 32'b1011001??????????000?????0110011
VFCPKD_S_S         = 32'b1011001??????????100?????0110011
VFCPKA_S_D         = 32'b1011010??????????000?????0110011
VFCPKB_S_D         = 32'b1011010??????????100?????0110011
VFCPKC_S_D         = 32'b1011011??????????000?????0110011
VFCPKD_S_D         = 32'b1011011??????????100?????0110011
VFADD_H            = 32'b1000001??????????010?????0110011
VFADD_R_H          = 32'b1000001??????????110?????0110011
VFSUB_H            = 32'b1000010??????????010?????0110011
VFSUB_R_H          = 32'b1000010??????????110?????0110011
VFMUL_H            = 32'b1000011??????????010?????0110011
VFMUL_R_H          = 32'b1000011??????????110?????0110011
VFDIV_H            = 32'b1000100??????????010?????0110011
VFDIV_R_H          = 32'b1000100??????????110?????0110011
VFMIN_H            = 32'b1000101??????????010?????0110011
VFMIN_R_H          = 32'b1000101??????????110?????0110011
VFMAX_H            = 32'b1000110??????????010?????0110011
VFMAX_R_H          = 32'b1000110??????????110?????0110011
VFSQRT_H           = 32'b100011100000?????010?????0110011
VFMAC_H            = 32'b1001000??????????010?????0110011
VFMAC_R_H          = 32'b1001000??????????110?????0110011
VFMRE_H            = 32'b1001001??????????010?????0110011
VFMRE_R_H          = 32'b1001001??????????110?????0110011
VFCLASS_H          = 32'b100110000001?????010?????0110011
VFSGNJ_H           = 32'b1001101??????????010?????0110011
VFSGNJ_R_H         = 32'b1001101??????????110?????0110011
VFSGNJN_H          = 32'b1001110??????????010?????0110011
VFSGNJN_R_H        = 32'b1001110??????????110?????0110011
VFSGNJX_H          = 32'b1001111??????????010?????0110011
VFSGNJX_R_H        = 32'b1001111??????????110?????0110011
VFEQ_H             = 32'b1010000??????????010?????0110011
VFEQ_R_H           = 32'b1010000??????????110?????0110011
VFNE_H             = 32'b1010001??????????010?????0110011
VFNE_R_H           = 32'b1010001??????????110?????0110011
VFLT_H             = 32'b1010010??????????010?????0110011
VFLT_R_H           = 32'b1010010??????????110?????0110011
VFGE_H             = 32'b1010011??????????010?????0110011
VFGE_R_H           = 32'b1010011??????????110?????0110011
VFLE_H             = 32'b1010100??????????010?????0110011
VFLE_R_H           = 32'b1010100??????????110?????0110011
VFGT_H             = 32'b1010101??????????010?????0110011
VFGT_R_H           = 32'b1010101??????????110?????0110011
VFMV_X_H           = 32'b100110000000?????010?????0110011
VFMV_H_X           = 32'b100110000000?????110?????0110011
VFCVT_X_H          = 32'b100110000010?????010?????0110011
VFCVT_XU_H         = 32'b100110000010?????110?????0110011
VFCVT_H_X          = 32'b100110000011?????010?????0110011
VFCVT_H_XU         = 32'b100110000011?????110?????0110011
VFCPKA_H_S         = 32'b1011000??????????010?????0110011
VFCPKB_H_S         = 32'b1011000??????????110?????0110011
VFCPKC_H_S         = 32'b1011001??????????010?????0110011
VFCPKD_H_S         = 32'b1011001??????????110?????0110011
VFCPKA_H_D         = 32'b1011010??????????010?????0110011
VFCPKB_H_D         = 32'b1011010??????????110?????0110011
VFCPKC_H_D         = 32'b1011011??????????010?????0110011
VFCPKD_H_D         = 32'b1011011??????????110?????0110011
VFCVT_S_H          = 32'b100110000110?????000?????0110011
VFCVTU_S_H         = 32'b100110000110?????100?????0110011
VFCVT_H_S          = 32'b100110000100?????010?????0110011
VFCVTU_H_S         = 32'b100110000100?????110?????0110011
VFADD_AH           = 32'b1000001??????????001?????0110011
VFADD_R_AH         = 32'b1000001??????????101?????0110011
VFSUB_AH           = 32'b1000010??????????001?????0110011
VFSUB_R_AH         = 32'b1000010??????????101?????0110011
VFMUL_AH           = 32'b1000011??????????001?????0110011
VFMUL_R_AH         = 32'b1000011??????????101?????0110011
VFDIV_AH           = 32'b1000100??????????001?????0110011
VFDIV_R_AH         = 32'b1000100??????????101?????0110011
VFMIN_AH           = 32'b1000101??????????001?????0110011
VFMIN_R_AH         = 32'b1000101??????????101?????0110011
VFMAX_AH           = 32'b1000110??????????001?????0110011
VFMAX_R_AH         = 32'b1000110??????????101?????0110011
VFSQRT_AH          = 32'b100011100000?????001?????0110011
VFMAC_AH           = 32'b1001000??????????001?????0110011
VFMAC_R_AH         = 32'b1001000??????????101?????0110011
VFMRE_AH           = 32'b1001001??????????001?????0110011
VFMRE_R_AH         = 32'b1001001??????????101?????0110011
VFCLASS_AH         = 32'b100110000001?????001?????0110011
VFSGNJ_AH          = 32'b1001101??????????001?????0110011
VFSGNJ_R_AH        = 32'b1001101??????????101?????0110011
VFSGNJN_AH         = 32'b1001110??????????001?????0110011
VFSGNJN_R_AH       = 32'b1001110??????????101?????0110011
VFSGNJX_AH         = 32'b1001111??????????001?????0110011
VFSGNJX_R_AH       = 32'b1001111??????????101?????0110011
VFEQ_AH            = 32'b1010000??????????001?????0110011
VFEQ_R_AH          = 32'b1010000??????????101?????0110011
VFNE_AH            = 32'b1010001??????????001?????0110011
VFNE_R_AH          = 32'b1010001??????????101?????0110011
VFLT_AH            = 32'b1010010??????????001?????0110011
VFLT_R_AH          = 32'b1010010??????????101?????0110011
VFGE_AH            = 32'b1010011??????????001?????0110011
VFGE_R_AH          = 32'b1010011??????????101?????0110011
VFLE_AH            = 32'b1010100??????????001?????0110011
VFLE_R_AH          = 32'b1010100??????????101?????0110011
VFGT_AH            = 32'b1010101??????????001?????0110011
VFGT_R_AH          = 32'b1010101??????????101?????0110011
VFMV_X_AH          = 32'b100110000000?????001?????0110011
VFMV_AH_X          = 32'b100110000000?????101?????0110011
VFCVT_X_AH         = 32'b100110000010?????001?????0110011
VFCVT_XU_AH        = 32'b100110000010?????101?????0110011
VFCVT_AH_X         = 32'b100110000011?????001?????0110011
VFCVT_AH_XU        = 32'b100110000011?????101?????0110011
VFCPKA_AH_S        = 32'b1011000??????????001?????0110011
VFCPKB_AH_S        = 32'b1011000??????????101?????0110011
VFCPKC_AH_S        = 32'b1011001??????????001?????0110011
VFCPKD_AH_S        = 32'b1011001??????????101?????0110011
VFCPKA_AH_D        = 32'b1011010??????????001?????0110011
VFCPKB_AH_D        = 32'b1011010??????????101?????0110011
VFCPKC_AH_D        = 32'b1011011??????????001?????0110011
VFCPKD_AH_D        = 32'b1011011??????????101?????0110011
VFCVT_S_AH         = 32'b100110000101?????000?????0110011
VFCVTU_S_AH        = 32'b100110000101?????100?????0110011
VFCVT_AH_S         = 32'b100110000100?????001?????0110011
VFCVTU_AH_S        = 32'b100110000100?????101?????0110011
VFCVT_H_AH         = 32'b100110000101?????010?????0110011
VFCVTU_H_AH        = 32'b100110000101?????110?????0110011
VFCVT_AH_H         = 32'b100110000110?????001?????0110011
VFCVTU_AH_H        = 32'b100110000110?????101?????0110011
VFADD_B            = 32'b1000001??????????011?????0110011
VFADD_R_B          = 32'b1000001??????????111?????0110011
VFSUB_B            = 32'b1000010??????????011?????0110011
VFSUB_R_B          = 32'b1000010??????????111?????0110011
VFMUL_B            = 32'b1000011??????????011?????0110011
VFMUL_R_B          = 32'b1000011??????????111?????0110011
VFDIV_B            = 32'b1000100??????????011?????0110011
VFDIV_R_B          = 32'b1000100??????????111?????0110011
VFMIN_B            = 32'b1000101??????????011?????0110011
VFMIN_R_B          = 32'b1000101??????????111?????0110011
VFMAX_B            = 32'b1000110??????????011?????0110011
VFMAX_R_B          = 32'b1000110??????????111?????0110011
VFSQRT_B           = 32'b100011100000?????011?????0110011
VFMAC_B            = 32'b1001000??????????011?????0110011
VFMAC_R_B          = 32'b1001000??????????111?????0110011
VFMRE_B            = 32'b1001001??????????011?????0110011
VFMRE_R_B          = 32'b1001001??????????111?????0110011
VFSGNJ_B           = 32'b1001101??????????011?????0110011
VFSGNJ_R_B         = 32'b1001101??????????111?????0110011
VFSGNJN_B          = 32'b1001110??????????011?????0110011
VFSGNJN_R_B        = 32'b1001110??????????111?????0110011
VFSGNJX_B          = 32'b1001111??????????011?????0110011
VFSGNJX_R_B        = 32'b1001111??????????111?????0110011
VFEQ_B             = 32'b1010000??????????011?????0110011
VFEQ_R_B           = 32'b1010000??????????111?????0110011
VFNE_B             = 32'b1010001??????????011?????0110011
VFNE_R_B           = 32'b1010001??????????111?????0110011
VFLT_B             = 32'b1010010??????????011?????0110011
VFLT_R_B           = 32'b1010010??????????111?????0110011
VFGE_B             = 32'b1010011??????????011?????0110011
VFGE_R_B           = 32'b1010011??????????111?????0110011
VFLE_B             = 32'b1010100??????????011?????0110011
VFLE_R_B           = 32'b1010100??????????111?????0110011
VFGT_B             = 32'b1010101??????????011?????0110011
VFGT_R_B           = 32'b1010101??????????111?????0110011
VFMV_X_B           = 32'b100110000000?????011?????0110011
VFMV_B_X           = 32'b100110000000?????111?????0110011
VFCLASS_B          = 32'b100110000001?????011?????0110011
VFCVT_X_B          = 32'b100110000010?????011?????0110011
VFCVT_XU_B         = 32'b100110000010?????111?????0110011
VFCVT_B_X          = 32'b100110000011?????011?????0110011
VFCVT_B_XU         = 32'b100110000011?????111?????0110011
VFCPKA_B_S         = 32'b1011000??????????011?????0110011
VFCPKB_B_S         = 32'b1011000??????????111?????0110011
VFCPKC_B_S         = 32'b1011001??????????011?????0110011
VFCPKD_B_S         = 32'b1011001??????????111?????0110011
VFCPKA_B_D         = 32'b1011010??????????011?????0110011
VFCPKB_B_D         = 32'b1011010??????????111?????0110011
VFCPKC_B_D         = 32'b1011011??????????011?????0110011
VFCPKD_B_D         = 32'b1011011??????????111?????0110011
VFCVT_S_B          = 32'b100110000111?????000?????0110011
VFCVTU_S_B         = 32'b100110000111?????100?????0110011
VFCVT_B_S          = 32'b100110000100?????011?????0110011
VFCVTU_B_S         = 32'b100110000100?????111?????0110011
VFCVT_H_B          = 32'b100110000111?????010?????0110011
VFCVTU_H_B         = 32'b100110000111?????110?????0110011
VFCVT_B_H          = 32'b100110000110?????011?????0110011
VFCVTU_B_H         = 32'b100110000110?????111?????0110011
VFCVT_AH_B         = 32'b100110000111?????001?????0110011
VFCVTU_AH_B        = 32'b100110000111?????101?????0110011
VFCVT_B_AH         = 32'b100110000101?????011?????0110011
VFCVTU_B_AH        = 32'b100110000101?????111?????0110011
VFDOTP_S           = 32'b1001010??????????000?????0110011
VFDOTP_R_S         = 32'b1001010??????????100?????0110011
VFAVG_S            = 32'b1010110??????????000?????0110011
VFAVG_R_S          = 32'b1010110??????????100?????0110011
FMULEX_S_H         = 32'b0100110??????????????????1010011
FMACEX_S_H         = 32'b0101010??????????????????1010011
VFDOTP_H           = 32'b1001010??????????010?????0110011
VFDOTP_R_H         = 32'b1001010??????????110?????0110011
VFDOTPEX_S_H       = 32'b1001011??????????010?????0110011
VFDOTPEX_S_R_H     = 32'b1001011??????????110?????0110011
VFAVG_H            = 32'b1010110??????????010?????0110011
VFAVG_R_H          = 32'b1010110??????????110?????0110011
FMULEX_S_AH        = 32'b0100110??????????101?????1010011
FMACEX_S_AH        = 32'b0101010??????????101?????1010011
VFDOTP_AH          = 32'b1001010??????????001?????0110011
VFDOTP_R_AH        = 32'b1001010??????????101?????0110011
VFDOTPEX_S_AH      = 32'b1001011??????????001?????0110011
VFDOTPEX_S_R_AH    = 32'b1001011??????????101?????0110011
VFAVG_AH           = 32'b1010110??????????001?????0110011
VFAVG_R_AH         = 32'b1010110??????????101?????0110011
FMULEX_S_B         = 32'b0100111??????????????????1010011
FMACEX_S_B         = 32'b0101011??????????????????1010011
VFDOTP_B           = 32'b1001010??????????011?????0110011
VFDOTP_R_B         = 32'b1001010??????????111?????0110011
VFDOTPEX_S_B       = 32'b1001011??????????011?????0110011
VFDOTPEX_S_R_B     = 32'b1001011??????????111?????0110011
VFAVG_B            = 32'b1010110??????????011?????0110011
VFAVG_R_B          = 32'b1010110??????????111?????0110011