package fpu_ss_instr_pkg;
  localparam logic [15:0] C_FLWSP            = 16'b011???????????10;
  localparam logic [15:0] C_FSWSP            = 16'b111???????????10;
  localparam logic [15:0] C_FLW              = 16'b011???????????00;
  localparam logic [15:0] C_FSW              = 16'b111???????????00;

  localparam logic [31:0] CSRRW_FSCSR        = 32'b000000000011?????001?????1110011;
  localparam logic [31:0] CSRRS_FRCSR        = 32'b000000000011?????010?????1110011;
  localparam logic [31:0] CSRRW_FSRM         = 32'b000000000010?????001?????1110011;
  localparam logic [31:0] CSRRS_FRRM         = 32'b000000000010?????010?????1110011;
  localparam logic [31:0] CSRRWI_FSRMI       = 32'b000000000010?????101?????1110011;
  localparam logic [31:0] CSRRW_FSFLAGS      = 32'b000000000001?????001?????1110011;
  localparam logic [31:0] CSRRS_FRFLAGS      = 32'b000000000001?????010?????1110011;
  localparam logic [31:0] CSRRWI_FSFLAGSI    = 32'b000000000001?????101?????1110011;
  localparam logic [31:0] FADD_S             = 32'b0000000??????????????????1010011;
  localparam logic [31:0] FSUB_S             = 32'b0000100??????????????????1010011;
  localparam logic [31:0] FMUL_S             = 32'b0001000??????????????????1010011;
  localparam logic [31:0] FDIV_S             = 32'b0001100??????????????????1010011;
  localparam logic [31:0] FSGNJ_S            = 32'b0010000??????????000?????1010011;
  localparam logic [31:0] FSGNJN_S           = 32'b0010000??????????001?????1010011;
  localparam logic [31:0] FSGNJX_S           = 32'b0010000??????????010?????1010011;
  localparam logic [31:0] FMIN_S             = 32'b0010100??????????000?????1010011;
  localparam logic [31:0] FMAX_S             = 32'b0010100??????????001?????1010011;
  localparam logic [31:0] FSQRT_S            = 32'b010110000000?????????????1010011;
  localparam logic [31:0] FADD_D             = 32'b0000001??????????????????1010011;
  localparam logic [31:0] FSUB_D             = 32'b0000101??????????????????1010011;
  localparam logic [31:0] FMUL_D             = 32'b0001001??????????????????1010011;
  localparam logic [31:0] FDIV_D             = 32'b0001101??????????????????1010011;
  localparam logic [31:0] FSGNJ_D            = 32'b0010001??????????000?????1010011;
  localparam logic [31:0] FSGNJN_D           = 32'b0010001??????????001?????1010011;
  localparam logic [31:0] FSGNJX_D           = 32'b0010001??????????010?????1010011;
  localparam logic [31:0] FMIN_D             = 32'b0010101??????????000?????1010011;
  localparam logic [31:0] FMAX_D             = 32'b0010101??????????001?????1010011;
  localparam logic [31:0] FCVT_S_D           = 32'b010000000001?????????????1010011;
  localparam logic [31:0] FCVT_D_S           = 32'b010000100000?????????????1010011;
  localparam logic [31:0] FSQRT_D            = 32'b010110100000?????????????1010011;
  localparam logic [31:0] FADD_Q             = 32'b0000011??????????????????1010011;
  localparam logic [31:0] FSUB_Q             = 32'b0000111??????????????????1010011;
  localparam logic [31:0] FMUL_Q             = 32'b0001011??????????????????1010011;
  localparam logic [31:0] FDIV_Q             = 32'b0001111??????????????????1010011;
  localparam logic [31:0] FSGNJ_Q            = 32'b0010011??????????000?????1010011;
  localparam logic [31:0] FSGNJN_Q           = 32'b0010011??????????001?????1010011;
  localparam logic [31:0] FSGNJX_Q           = 32'b0010011??????????010?????1010011;
  localparam logic [31:0] FMIN_Q             = 32'b0010111??????????000?????1010011;
  localparam logic [31:0] FMAX_Q             = 32'b0010111??????????001?????1010011;
  localparam logic [31:0] FCVT_S_Q           = 32'b010000000011?????????????1010011;
  localparam logic [31:0] FCVT_Q_S           = 32'b010001100000?????????????1010011;
  localparam logic [31:0] FCVT_D_Q           = 32'b010000100011?????????????1010011;
  localparam logic [31:0] FCVT_Q_D           = 32'b010001100001?????????????1010011;
  localparam logic [31:0] FSQRT_Q            = 32'b010111100000?????????????1010011;
  localparam logic [31:0] FLE_S              = 32'b1010000??????????000?????1010011;
  localparam logic [31:0] FLT_S              = 32'b1010000??????????001?????1010011;
  localparam logic [31:0] FEQ_S              = 32'b1010000??????????010?????1010011;
  localparam logic [31:0] FLE_D              = 32'b1010001??????????000?????1010011;
  localparam logic [31:0] FLT_D              = 32'b1010001??????????001?????1010011;
  localparam logic [31:0] FEQ_D              = 32'b1010001??????????010?????1010011;
  localparam logic [31:0] FLE_Q              = 32'b1010011??????????000?????1010011;
  localparam logic [31:0] FLT_Q              = 32'b1010011??????????001?????1010011;
  localparam logic [31:0] FEQ_Q              = 32'b1010011??????????010?????1010011;
  localparam logic [31:0] FCVT_W_S           = 32'b110000000000?????????????1010011;
  localparam logic [31:0] FCVT_WU_S          = 32'b110000000001?????????????1010011;
  localparam logic [31:0] FCVT_L_S           = 32'b110000000010?????????????1010011;
  localparam logic [31:0] FCVT_LU_S          = 32'b110000000011?????????????1010011;
  localparam logic [31:0] FMV_X_W            = 32'b111000000000?????000?????1010011;
  localparam logic [31:0] FCLASS_S           = 32'b111000000000?????001?????1010011;
  localparam logic [31:0] FCVT_W_D           = 32'b110000100000?????????????1010011;
  localparam logic [31:0] FCVT_WU_D          = 32'b110000100001?????????????1010011;
  localparam logic [31:0] FCVT_L_D           = 32'b110000100010?????????????1010011;
  localparam logic [31:0] FCVT_LU_D          = 32'b110000100011?????????????1010011;
  localparam logic [31:0] FMV_X_D            = 32'b111000100000?????000?????1010011;
  localparam logic [31:0] FCLASS_D           = 32'b111000100000?????001?????1010011;
  localparam logic [31:0] FCVT_W_Q           = 32'b110001100000?????????????1010011;
  localparam logic [31:0] FCVT_WU_Q          = 32'b110001100001?????????????1010011;
  localparam logic [31:0] FCVT_L_Q           = 32'b110001100010?????????????1010011;
  localparam logic [31:0] FCVT_LU_Q          = 32'b110001100011?????????????1010011;
  localparam logic [31:0] FMV_X_Q            = 32'b111001100000?????000?????1010011;
  localparam logic [31:0] FCLASS_Q           = 32'b111001100000?????001?????1010011;
  localparam logic [31:0] FCVT_S_W           = 32'b110100000000?????????????1010011;
  localparam logic [31:0] FCVT_S_WU          = 32'b110100000001?????????????1010011;
  localparam logic [31:0] FCVT_S_L           = 32'b110100000010?????????????1010011;
  localparam logic [31:0] FCVT_S_LU          = 32'b110100000011?????????????1010011;
  localparam logic [31:0] FMV_W_X            = 32'b111100000000?????000?????1010011;
  localparam logic [31:0] FCVT_D_W           = 32'b110100100000?????????????1010011;
  localparam logic [31:0] FCVT_D_WU          = 32'b110100100001?????????????1010011;
  localparam logic [31:0] FCVT_D_L           = 32'b110100100010?????????????1010011;
  localparam logic [31:0] FCVT_D_LU          = 32'b110100100011?????????????1010011;
  localparam logic [31:0] FMV_D_X            = 32'b111100100000?????000?????1010011;
  localparam logic [31:0] FCVT_Q_W           = 32'b110101100000?????????????1010011;
  localparam logic [31:0] FCVT_Q_WU          = 32'b110101100001?????????????1010011;
  localparam logic [31:0] FCVT_Q_L           = 32'b110101100010?????????????1010011;
  localparam logic [31:0] FCVT_Q_LU          = 32'b110101100011?????????????1010011;
  localparam logic [31:0] FMV_Q_X            = 32'b111101100000?????000?????1010011;
  localparam logic [31:0] FLW                = 32'b?????????????????010?????0000111;
  localparam logic [31:0] FLD                = 32'b?????????????????011?????0000111;
  localparam logic [31:0] FLQ                = 32'b?????????????????100?????0000111;
  localparam logic [31:0] FSW                = 32'b?????????????????010?????0100111;
  localparam logic [31:0] FSD                = 32'b?????????????????011?????0100111;
  localparam logic [31:0] FSQ                = 32'b?????????????????100?????0100111;
  localparam logic [31:0] FMADD_S            = 32'b?????00??????????????????1000011;
  localparam logic [31:0] FMSUB_S            = 32'b?????00??????????????????1000111;
  localparam logic [31:0] FNMSUB_S           = 32'b?????00??????????????????1001011;
  localparam logic [31:0] FNMADD_S           = 32'b?????00??????????????????1001111;
  localparam logic [31:0] FMADD_D            = 32'b?????01??????????????????1000011;
  localparam logic [31:0] FMSUB_D            = 32'b?????01??????????????????1000111;
  localparam logic [31:0] FNMSUB_D           = 32'b?????01??????????????????1001011;
  localparam logic [31:0] FNMADD_D           = 32'b?????01??????????????????1001111;
  localparam logic [31:0] FMADD_Q            = 32'b?????11??????????????????1000011;
  localparam logic [31:0] FMSUB_Q            = 32'b?????11??????????????????1000111;
  localparam logic [31:0] FNMSUB_Q           = 32'b?????11??????????????????1001011;
  localparam logic [31:0] FNMADD_Q           = 32'b?????11??????????????????1001111;
  localparam logic [31:0] DMSRC              = 32'b0000000??????????000000000101011;
  localparam logic [31:0] DMDST              = 32'b0000001??????????000000000101011;
  localparam logic [31:0] DMCPYI             = 32'b0000010??????????000?????0101011;
  localparam logic [31:0] DMCPY              = 32'b0000011??????????000?????0101011;
  localparam logic [31:0] DMSTATI            = 32'b0000100?????00000000?????0101011;
  localparam logic [31:0] DMSTAT             = 32'b0000101?????00000000?????0101011;
  localparam logic [31:0] DMSTR              = 32'b0000110??????????000000000101011;
  localparam logic [31:0] DMREP              = 32'b000011100000?????000000000101011;
  localparam logic [31:0] FREP_O             = 32'b????????????????????????10001011;
  localparam logic [31:0] FREP_I             = 32'b????????????????????????00001011;
  localparam logic [31:0] IREP               = 32'b?????????????????????????0111111;
  localparam logic [31:0] SCFGRI             = 32'b????????????00000001?????0101011;
  localparam logic [31:0] SCFGWI             = 32'b?????????????????010000000101011;
  localparam logic [31:0] SCFGR              = 32'b0000000?????00001001?????0101011;
  localparam logic [31:0] SCFGW              = 32'b0000000??????????010000010101011;
  localparam logic [31:0] FLH                = 32'b?????????????????001?????0000111;
  localparam logic [31:0] FSH                = 32'b?????????????????001?????0100111;
  localparam logic [31:0] FMADD_H            = 32'b?????10??????????????????1000011;
  localparam logic [31:0] FMSUB_H            = 32'b?????10??????????????????1000111;
  localparam logic [31:0] FNMSUB_H           = 32'b?????10??????????????????1001011;
  localparam logic [31:0] FNMADD_H           = 32'b?????10??????????????????1001111;
  localparam logic [31:0] FADD_H             = 32'b0000010??????????????????1010011;
  localparam logic [31:0] FSUB_H             = 32'b0000110??????????????????1010011;
  localparam logic [31:0] FMUL_H             = 32'b0001010??????????????????1010011;
  localparam logic [31:0] FDIV_H             = 32'b0001110??????????????????1010011;
  localparam logic [31:0] FSQRT_H            = 32'b010111000000?????????????1010011;
  localparam logic [31:0] FSGNJ_H            = 32'b0010010??????????000?????1010011;
  localparam logic [31:0] FSGNJN_H           = 32'b0010010??????????001?????1010011;
  localparam logic [31:0] FSGNJX_H           = 32'b0010010??????????010?????1010011;
  localparam logic [31:0] FMIN_H             = 32'b0010110??????????000?????1010011;
  localparam logic [31:0] FMAX_H             = 32'b0010110??????????001?????1010011;
  localparam logic [31:0] FEQ_H              = 32'b1010010??????????010?????1010011;
  localparam logic [31:0] FLT_H              = 32'b1010010??????????001?????1010011;
  localparam logic [31:0] FLE_H              = 32'b1010010??????????000?????1010011;
  localparam logic [31:0] FCVT_W_H           = 32'b110001000000?????????????1010011;
  localparam logic [31:0] FCVT_WU_H          = 32'b110001000001?????????????1010011;
  localparam logic [31:0] FCVT_H_W           = 32'b110101000000?????????????1010011;
  localparam logic [31:0] FCVT_H_WU          = 32'b110101000001?????????????1010011;
  localparam logic [31:0] FMV_X_H            = 32'b111001000000?????000?????1010011;
  localparam logic [31:0] FCLASS_H           = 32'b111001000000?????001?????1010011;
  localparam logic [31:0] FMV_H_X            = 32'b111101000000?????000?????1010011;
  localparam logic [31:0] FCVT_L_H           = 32'b110001000010?????????????1010011;
  localparam logic [31:0] FCVT_LU_H          = 32'b110001000011?????????????1010011;
  localparam logic [31:0] FCVT_H_L           = 32'b110101000010?????????????1010011;
  localparam logic [31:0] FCVT_H_LU          = 32'b110101000011?????????????1010011;
  localparam logic [31:0] FCVT_S_H           = 32'b010000000010?????000?????1010011;
  localparam logic [31:0] FCVT_H_S           = 32'b010001000000?????????????1010011;
  localparam logic [31:0] FCVT_D_H           = 32'b010000100010?????000?????1010011;
  localparam logic [31:0] FCVT_H_D           = 32'b010001000001?????????????1010011;
  localparam logic [31:0] FLAH               = 32'b?????????????????001?????0000111;
  localparam logic [31:0] FSAH               = 32'b?????????????????001?????0100111;
  localparam logic [31:0] FMADD_AH           = 32'b?????10??????????101?????1000011;
  localparam logic [31:0] FMSUB_AH           = 32'b?????10??????????101?????1000111;
  localparam logic [31:0] FNMSUB_AH          = 32'b?????10??????????101?????1001011;
  localparam logic [31:0] FNMADD_AH          = 32'b?????10??????????101?????1001111;
  localparam logic [31:0] FADD_AH            = 32'b0000010??????????101?????1010011;
  localparam logic [31:0] FSUB_AH            = 32'b0000110??????????101?????1010011;
  localparam logic [31:0] FMUL_AH            = 32'b0001010??????????101?????1010011;
  localparam logic [31:0] FDIV_AH            = 32'b0001110??????????101?????1010011;
  localparam logic [31:0] FSQRT_AH           = 32'b010111000000?????101?????1010011;
  localparam logic [31:0] FSGNJ_AH           = 32'b0010010??????????100?????1010011;
  localparam logic [31:0] FSGNJN_AH          = 32'b0010010??????????101?????1010011;
  localparam logic [31:0] FSGNJX_AH          = 32'b0010010??????????110?????1010011;
  localparam logic [31:0] FMIN_AH            = 32'b0010110??????????100?????1010011;
  localparam logic [31:0] FMAX_AH            = 32'b0010110??????????101?????1010011;
  localparam logic [31:0] FEQ_AH             = 32'b1010010??????????110?????1010011;
  localparam logic [31:0] FLT_AH             = 32'b1010010??????????101?????1010011;
  localparam logic [31:0] FLE_AH             = 32'b1010010??????????100?????1010011;
  localparam logic [31:0] FCVT_W_AH          = 32'b110001000000?????101?????1010011;
  localparam logic [31:0] FCVT_WU_AH         = 32'b110001000001?????101?????1010011;
  localparam logic [31:0] FCVT_AH_W          = 32'b110101000000?????101?????1010011;
  localparam logic [31:0] FCVT_AH_WU         = 32'b110101000001?????101?????1010011;
  localparam logic [31:0] FMV_X_AH           = 32'b111001000000?????100?????1010011;
  localparam logic [31:0] FCLASS_AH          = 32'b111001000000?????101?????1010011;
  localparam logic [31:0] FMV_AH_X           = 32'b111101000000?????100?????1010011;
  localparam logic [31:0] FCVT_L_AH          = 32'b110001000010?????101?????1010011;
  localparam logic [31:0] FCVT_LU_AH         = 32'b110001000011?????101?????1010011;
  localparam logic [31:0] FCVT_AH_L          = 32'b110101000010?????101?????1010011;
  localparam logic [31:0] FCVT_AH_LU         = 32'b110101000011?????101?????1010011;
  localparam logic [31:0] FCVT_S_AH          = 32'b010000000110?????000?????1010011;
  localparam logic [31:0] FCVT_AH_S          = 32'b010001000000?????101?????1010011;
  localparam logic [31:0] FCVT_D_AH          = 32'b010000100110?????000?????1010011;
  localparam logic [31:0] FCVT_AH_D          = 32'b010001000001?????101?????1010011;
  localparam logic [31:0] FCVT_H_AH          = 32'b010001000110?????????????1010011;
  localparam logic [31:0] FCVT_AH_H          = 32'b010001000010?????101?????1010011;
  localparam logic [31:0] FLB                = 32'b?????????????????000?????0000111;
  localparam logic [31:0] FSB                = 32'b?????????????????000?????0100111;
  localparam logic [31:0] FMADD_B            = 32'b?????11??????????????????1000011;
  localparam logic [31:0] FMSUB_B            = 32'b?????11??????????????????1000111;
  localparam logic [31:0] FNMSUB_B           = 32'b?????11??????????????????1001011;
  localparam logic [31:0] FNMADD_B           = 32'b?????11??????????????????1001111;
  localparam logic [31:0] FADD_B             = 32'b0000011??????????????????1010011;
  localparam logic [31:0] FSUB_B             = 32'b0000111??????????????????1010011;
  localparam logic [31:0] FMUL_B             = 32'b0001011??????????????????1010011;
  localparam logic [31:0] FDIV_B             = 32'b0001111??????????????????1010011;
  localparam logic [31:0] FSQRT_B            = 32'b010111100000?????????????1010011;
  localparam logic [31:0] FSGNJ_B            = 32'b0010011??????????000?????1010011;
  localparam logic [31:0] FSGNJN_B           = 32'b0010011??????????001?????1010011;
  localparam logic [31:0] FSGNJX_B           = 32'b0010011??????????010?????1010011;
  localparam logic [31:0] FMIN_B             = 32'b0010111??????????000?????1010011;
  localparam logic [31:0] FMAX_B             = 32'b0010111??????????001?????1010011;
  localparam logic [31:0] FEQ_B              = 32'b1010011??????????010?????1010011;
  localparam logic [31:0] FLT_B              = 32'b1010011??????????001?????1010011;
  localparam logic [31:0] FLE_B              = 32'b1010011??????????000?????1010011;
  localparam logic [31:0] FCVT_W_B           = 32'b110001100000?????????????1010011;
  localparam logic [31:0] FCVT_WU_B          = 32'b110001100001?????????????1010011;
  localparam logic [31:0] FCVT_B_W           = 32'b110101100000?????????????1010011;
  localparam logic [31:0] FCVT_B_WU          = 32'b110101100001?????????????1010011;
  localparam logic [31:0] FMV_X_B            = 32'b111001100000?????000?????1010011;
  localparam logic [31:0] FCLASS_B           = 32'b111001100000?????001?????1010011;
  localparam logic [31:0] FMV_B_X            = 32'b111101100000?????000?????1010011;
  localparam logic [31:0] FCVT_L_B           = 32'b110001100010?????????????1010011;
  localparam logic [31:0] FCVT_LU_B          = 32'b110001100011?????????????1010011;
  localparam logic [31:0] FCVT_B_L           = 32'b110101100010?????????????1010011;
  localparam logic [31:0] FCVT_B_LU          = 32'b110101100011?????????????1010011;
  localparam logic [31:0] FCVT_S_B           = 32'b010000000011?????000?????1010011;
  localparam logic [31:0] FCVT_B_S           = 32'b010001100000?????????????1010011;
  localparam logic [31:0] FCVT_D_B           = 32'b010000100011?????000?????1010011;
  localparam logic [31:0] FCVT_B_D           = 32'b010001100001?????????????1010011;
  localparam logic [31:0] FCVT_H_B           = 32'b010001000011?????000?????1010011;
  localparam logic [31:0] FCVT_B_H           = 32'b010001100010?????????????1010011;
  localparam logic [31:0] FCVT_AH_B          = 32'b010001000011?????101?????1010011;
  localparam logic [31:0] FCVT_B_AH          = 32'b010001100110?????????????1010011;
  localparam logic [31:0] VFADD_S            = 32'b1000001??????????000?????0110011;
  localparam logic [31:0] VFADD_R_S          = 32'b1000001??????????100?????0110011;
  localparam logic [31:0] VFSUB_S            = 32'b1000010??????????000?????0110011;
  localparam logic [31:0] VFSUB_R_S          = 32'b1000010??????????100?????0110011;
  localparam logic [31:0] VFMUL_S            = 32'b1000011??????????000?????0110011;
  localparam logic [31:0] VFMUL_R_S          = 32'b1000011??????????100?????0110011;
  localparam logic [31:0] VFDIV_S            = 32'b1000100??????????000?????0110011;
  localparam logic [31:0] VFDIV_R_S          = 32'b1000100??????????100?????0110011;
  localparam logic [31:0] VFMIN_S            = 32'b1000101??????????000?????0110011;
  localparam logic [31:0] VFMIN_R_S          = 32'b1000101??????????100?????0110011;
  localparam logic [31:0] VFMAX_S            = 32'b1000110??????????000?????0110011;
  localparam logic [31:0] VFMAX_R_S          = 32'b1000110??????????100?????0110011;
  localparam logic [31:0] VFSQRT_S           = 32'b100011100000?????000?????0110011;
  localparam logic [31:0] VFMAC_S            = 32'b1001000??????????000?????0110011;
  localparam logic [31:0] VFMAC_R_S          = 32'b1001000??????????100?????0110011;
  localparam logic [31:0] VFMRE_S            = 32'b1001001??????????000?????0110011;
  localparam logic [31:0] VFMRE_R_S          = 32'b1001001??????????100?????0110011;
  localparam logic [31:0] VFCLASS_S          = 32'b100110000001?????000?????0110011;
  localparam logic [31:0] VFSGNJ_S           = 32'b1001101??????????000?????0110011;
  localparam logic [31:0] VFSGNJ_R_S         = 32'b1001101??????????100?????0110011;
  localparam logic [31:0] VFSGNJN_S          = 32'b1001110??????????000?????0110011;
  localparam logic [31:0] VFSGNJN_R_S        = 32'b1001110??????????100?????0110011;
  localparam logic [31:0] VFSGNJX_S          = 32'b1001111??????????000?????0110011;
  localparam logic [31:0] VFSGNJX_R_S        = 32'b1001111??????????100?????0110011;
  localparam logic [31:0] VFEQ_S             = 32'b1010000??????????000?????0110011;
  localparam logic [31:0] VFEQ_R_S           = 32'b1010000??????????100?????0110011;
  localparam logic [31:0] VFNE_S             = 32'b1010001??????????000?????0110011;
  localparam logic [31:0] VFNE_R_S           = 32'b1010001??????????100?????0110011;
  localparam logic [31:0] VFLT_S             = 32'b1010010??????????000?????0110011;
  localparam logic [31:0] VFLT_R_S           = 32'b1010010??????????100?????0110011;
  localparam logic [31:0] VFGE_S             = 32'b1010011??????????000?????0110011;
  localparam logic [31:0] VFGE_R_S           = 32'b1010011??????????100?????0110011;
  localparam logic [31:0] VFLE_S             = 32'b1010100??????????000?????0110011;
  localparam logic [31:0] VFLE_R_S           = 32'b1010100??????????100?????0110011;
  localparam logic [31:0] VFGT_S             = 32'b1010101??????????000?????0110011;
  localparam logic [31:0] VFGT_R_S           = 32'b1010101??????????100?????0110011;
  localparam logic [31:0] VFMV_X_S           = 32'b100110000000?????000?????0110011;
  localparam logic [31:0] VFMV_S_X           = 32'b100110000000?????100?????0110011;
  localparam logic [31:0] VFCVT_X_S          = 32'b100110000010?????000?????0110011;
  localparam logic [31:0] VFCVT_XU_S         = 32'b100110000010?????100?????0110011;
  localparam logic [31:0] VFCVT_S_X          = 32'b100110000011?????000?????0110011;
  localparam logic [31:0] VFCVT_S_XU         = 32'b100110000011?????100?????0110011;
  localparam logic [31:0] VFCPKA_S_S         = 32'b1011000??????????000?????0110011;
  localparam logic [31:0] VFCPKB_S_S         = 32'b1011000??????????100?????0110011;
  localparam logic [31:0] VFCPKC_S_S         = 32'b1011001??????????000?????0110011;
  localparam logic [31:0] VFCPKD_S_S         = 32'b1011001??????????100?????0110011;
  localparam logic [31:0] VFCPKA_S_D         = 32'b1011010??????????000?????0110011;
  localparam logic [31:0] VFCPKB_S_D         = 32'b1011010??????????100?????0110011;
  localparam logic [31:0] VFCPKC_S_D         = 32'b1011011??????????000?????0110011;
  localparam logic [31:0] VFCPKD_S_D         = 32'b1011011??????????100?????0110011;
  localparam logic [31:0] VFADD_H            = 32'b1000001??????????010?????0110011;
  localparam logic [31:0] VFADD_R_H          = 32'b1000001??????????110?????0110011;
  localparam logic [31:0] VFSUB_H            = 32'b1000010??????????010?????0110011;
  localparam logic [31:0] VFSUB_R_H          = 32'b1000010??????????110?????0110011;
  localparam logic [31:0] VFMUL_H            = 32'b1000011??????????010?????0110011;
  localparam logic [31:0] VFMUL_R_H          = 32'b1000011??????????110?????0110011;
  localparam logic [31:0] VFDIV_H            = 32'b1000100??????????010?????0110011;
  localparam logic [31:0] VFDIV_R_H          = 32'b1000100??????????110?????0110011;
  localparam logic [31:0] VFMIN_H            = 32'b1000101??????????010?????0110011;
  localparam logic [31:0] VFMIN_R_H          = 32'b1000101??????????110?????0110011;
  localparam logic [31:0] VFMAX_H            = 32'b1000110??????????010?????0110011;
  localparam logic [31:0] VFMAX_R_H          = 32'b1000110??????????110?????0110011;
  localparam logic [31:0] VFSQRT_H           = 32'b100011100000?????010?????0110011;
  localparam logic [31:0] VFMAC_H            = 32'b1001000??????????010?????0110011;
  localparam logic [31:0] VFMAC_R_H          = 32'b1001000??????????110?????0110011;
  localparam logic [31:0] VFMRE_H            = 32'b1001001??????????010?????0110011;
  localparam logic [31:0] VFMRE_R_H          = 32'b1001001??????????110?????0110011;
  localparam logic [31:0] VFCLASS_H          = 32'b100110000001?????010?????0110011;
  localparam logic [31:0] VFSGNJ_H           = 32'b1001101??????????010?????0110011;
  localparam logic [31:0] VFSGNJ_R_H         = 32'b1001101??????????110?????0110011;
  localparam logic [31:0] VFSGNJN_H          = 32'b1001110??????????010?????0110011;
  localparam logic [31:0] VFSGNJN_R_H        = 32'b1001110??????????110?????0110011;
  localparam logic [31:0] VFSGNJX_H          = 32'b1001111??????????010?????0110011;
  localparam logic [31:0] VFSGNJX_R_H        = 32'b1001111??????????110?????0110011;
  localparam logic [31:0] VFEQ_H             = 32'b1010000??????????010?????0110011;
  localparam logic [31:0] VFEQ_R_H           = 32'b1010000??????????110?????0110011;
  localparam logic [31:0] VFNE_H             = 32'b1010001??????????010?????0110011;
  localparam logic [31:0] VFNE_R_H           = 32'b1010001??????????110?????0110011;
  localparam logic [31:0] VFLT_H             = 32'b1010010??????????010?????0110011;
  localparam logic [31:0] VFLT_R_H           = 32'b1010010??????????110?????0110011;
  localparam logic [31:0] VFGE_H             = 32'b1010011??????????010?????0110011;
  localparam logic [31:0] VFGE_R_H           = 32'b1010011??????????110?????0110011;
  localparam logic [31:0] VFLE_H             = 32'b1010100??????????010?????0110011;
  localparam logic [31:0] VFLE_R_H           = 32'b1010100??????????110?????0110011;
  localparam logic [31:0] VFGT_H             = 32'b1010101??????????010?????0110011;
  localparam logic [31:0] VFGT_R_H           = 32'b1010101??????????110?????0110011;
  localparam logic [31:0] VFMV_X_H           = 32'b100110000000?????010?????0110011;
  localparam logic [31:0] VFMV_H_X           = 32'b100110000000?????110?????0110011;
  localparam logic [31:0] VFCVT_X_H          = 32'b100110000010?????010?????0110011;
  localparam logic [31:0] VFCVT_XU_H         = 32'b100110000010?????110?????0110011;
  localparam logic [31:0] VFCVT_H_X          = 32'b100110000011?????010?????0110011;
  localparam logic [31:0] VFCVT_H_XU         = 32'b100110000011?????110?????0110011;
  localparam logic [31:0] VFCPKA_H_S         = 32'b1011000??????????010?????0110011;
  localparam logic [31:0] VFCPKB_H_S         = 32'b1011000??????????110?????0110011;
  localparam logic [31:0] VFCPKC_H_S         = 32'b1011001??????????010?????0110011;
  localparam logic [31:0] VFCPKD_H_S         = 32'b1011001??????????110?????0110011;
  localparam logic [31:0] VFCPKA_H_D         = 32'b1011010??????????010?????0110011;
  localparam logic [31:0] VFCPKB_H_D         = 32'b1011010??????????110?????0110011;
  localparam logic [31:0] VFCPKC_H_D         = 32'b1011011??????????010?????0110011;
  localparam logic [31:0] VFCPKD_H_D         = 32'b1011011??????????110?????0110011;
  localparam logic [31:0] VFCVT_S_H          = 32'b100110000110?????000?????0110011;
  localparam logic [31:0] VFCVTU_S_H         = 32'b100110000110?????100?????0110011;
  localparam logic [31:0] VFCVT_H_S          = 32'b100110000100?????010?????0110011;
  localparam logic [31:0] VFCVTU_H_S         = 32'b100110000100?????110?????0110011;
  localparam logic [31:0] VFADD_AH           = 32'b1000001??????????001?????0110011;
  localparam logic [31:0] VFADD_R_AH         = 32'b1000001??????????101?????0110011;
  localparam logic [31:0] VFSUB_AH           = 32'b1000010??????????001?????0110011;
  localparam logic [31:0] VFSUB_R_AH         = 32'b1000010??????????101?????0110011;
  localparam logic [31:0] VFMUL_AH           = 32'b1000011??????????001?????0110011;
  localparam logic [31:0] VFMUL_R_AH         = 32'b1000011??????????101?????0110011;
  localparam logic [31:0] VFDIV_AH           = 32'b1000100??????????001?????0110011;
  localparam logic [31:0] VFDIV_R_AH         = 32'b1000100??????????101?????0110011;
  localparam logic [31:0] VFMIN_AH           = 32'b1000101??????????001?????0110011;
  localparam logic [31:0] VFMIN_R_AH         = 32'b1000101??????????101?????0110011;
  localparam logic [31:0] VFMAX_AH           = 32'b1000110??????????001?????0110011;
  localparam logic [31:0] VFMAX_R_AH         = 32'b1000110??????????101?????0110011;
  localparam logic [31:0] VFSQRT_AH          = 32'b100011100000?????001?????0110011;
  localparam logic [31:0] VFMAC_AH           = 32'b1001000??????????001?????0110011;
  localparam logic [31:0] VFMAC_R_AH         = 32'b1001000??????????101?????0110011;
  localparam logic [31:0] VFMRE_AH           = 32'b1001001??????????001?????0110011;
  localparam logic [31:0] VFMRE_R_AH         = 32'b1001001??????????101?????0110011;
  localparam logic [31:0] VFCLASS_AH         = 32'b100110000001?????001?????0110011;
  localparam logic [31:0] VFSGNJ_AH          = 32'b1001101??????????001?????0110011;
  localparam logic [31:0] VFSGNJ_R_AH        = 32'b1001101??????????101?????0110011;
  localparam logic [31:0] VFSGNJN_AH         = 32'b1001110??????????001?????0110011;
  localparam logic [31:0] VFSGNJN_R_AH       = 32'b1001110??????????101?????0110011;
  localparam logic [31:0] VFSGNJX_AH         = 32'b1001111??????????001?????0110011;
  localparam logic [31:0] VFSGNJX_R_AH       = 32'b1001111??????????101?????0110011;
  localparam logic [31:0] VFEQ_AH            = 32'b1010000??????????001?????0110011;
  localparam logic [31:0] VFEQ_R_AH          = 32'b1010000??????????101?????0110011;
  localparam logic [31:0] VFNE_AH            = 32'b1010001??????????001?????0110011;
  localparam logic [31:0] VFNE_R_AH          = 32'b1010001??????????101?????0110011;
  localparam logic [31:0] VFLT_AH            = 32'b1010010??????????001?????0110011;
  localparam logic [31:0] VFLT_R_AH          = 32'b1010010??????????101?????0110011;
  localparam logic [31:0] VFGE_AH            = 32'b1010011??????????001?????0110011;
  localparam logic [31:0] VFGE_R_AH          = 32'b1010011??????????101?????0110011;
  localparam logic [31:0] VFLE_AH            = 32'b1010100??????????001?????0110011;
  localparam logic [31:0] VFLE_R_AH          = 32'b1010100??????????101?????0110011;
  localparam logic [31:0] VFGT_AH            = 32'b1010101??????????001?????0110011;
  localparam logic [31:0] VFGT_R_AH          = 32'b1010101??????????101?????0110011;
  localparam logic [31:0] VFMV_X_AH          = 32'b100110000000?????001?????0110011;
  localparam logic [31:0] VFMV_AH_X          = 32'b100110000000?????101?????0110011;
  localparam logic [31:0] VFCVT_X_AH         = 32'b100110000010?????001?????0110011;
  localparam logic [31:0] VFCVT_XU_AH        = 32'b100110000010?????101?????0110011;
  localparam logic [31:0] VFCVT_AH_X         = 32'b100110000011?????001?????0110011;
  localparam logic [31:0] VFCVT_AH_XU        = 32'b100110000011?????101?????0110011;
  localparam logic [31:0] VFCPKA_AH_S        = 32'b1011000??????????001?????0110011;
  localparam logic [31:0] VFCPKB_AH_S        = 32'b1011000??????????101?????0110011;
  localparam logic [31:0] VFCPKC_AH_S        = 32'b1011001??????????001?????0110011;
  localparam logic [31:0] VFCPKD_AH_S        = 32'b1011001??????????101?????0110011;
  localparam logic [31:0] VFCPKA_AH_D        = 32'b1011010??????????001?????0110011;
  localparam logic [31:0] VFCPKB_AH_D        = 32'b1011010??????????101?????0110011;
  localparam logic [31:0] VFCPKC_AH_D        = 32'b1011011??????????001?????0110011;
  localparam logic [31:0] VFCPKD_AH_D        = 32'b1011011??????????101?????0110011;
  localparam logic [31:0] VFCVT_S_AH         = 32'b100110000101?????000?????0110011;
  localparam logic [31:0] VFCVTU_S_AH        = 32'b100110000101?????100?????0110011;
  localparam logic [31:0] VFCVT_AH_S         = 32'b100110000100?????001?????0110011;
  localparam logic [31:0] VFCVTU_AH_S        = 32'b100110000100?????101?????0110011;
  localparam logic [31:0] VFCVT_H_AH         = 32'b100110000101?????010?????0110011;
  localparam logic [31:0] VFCVTU_H_AH        = 32'b100110000101?????110?????0110011;
  localparam logic [31:0] VFCVT_AH_H         = 32'b100110000110?????001?????0110011;
  localparam logic [31:0] VFCVTU_AH_H        = 32'b100110000110?????101?????0110011;
  localparam logic [31:0] VFADD_B            = 32'b1000001??????????011?????0110011;
  localparam logic [31:0] VFADD_R_B          = 32'b1000001??????????111?????0110011;
  localparam logic [31:0] VFSUB_B            = 32'b1000010??????????011?????0110011;
  localparam logic [31:0] VFSUB_R_B          = 32'b1000010??????????111?????0110011;
  localparam logic [31:0] VFMUL_B            = 32'b1000011??????????011?????0110011;
  localparam logic [31:0] VFMUL_R_B          = 32'b1000011??????????111?????0110011;
  localparam logic [31:0] VFDIV_B            = 32'b1000100??????????011?????0110011;
  localparam logic [31:0] VFDIV_R_B          = 32'b1000100??????????111?????0110011;
  localparam logic [31:0] VFMIN_B            = 32'b1000101??????????011?????0110011;
  localparam logic [31:0] VFMIN_R_B          = 32'b1000101??????????111?????0110011;
  localparam logic [31:0] VFMAX_B            = 32'b1000110??????????011?????0110011;
  localparam logic [31:0] VFMAX_R_B          = 32'b1000110??????????111?????0110011;
  localparam logic [31:0] VFSQRT_B           = 32'b100011100000?????011?????0110011;
  localparam logic [31:0] VFMAC_B            = 32'b1001000??????????011?????0110011;
  localparam logic [31:0] VFMAC_R_B          = 32'b1001000??????????111?????0110011;
  localparam logic [31:0] VFMRE_B            = 32'b1001001??????????011?????0110011;
  localparam logic [31:0] VFMRE_R_B          = 32'b1001001??????????111?????0110011;
  localparam logic [31:0] VFSGNJ_B           = 32'b1001101??????????011?????0110011;
  localparam logic [31:0] VFSGNJ_R_B         = 32'b1001101??????????111?????0110011;
  localparam logic [31:0] VFSGNJN_B          = 32'b1001110??????????011?????0110011;
  localparam logic [31:0] VFSGNJN_R_B        = 32'b1001110??????????111?????0110011;
  localparam logic [31:0] VFSGNJX_B          = 32'b1001111??????????011?????0110011;
  localparam logic [31:0] VFSGNJX_R_B        = 32'b1001111??????????111?????0110011;
  localparam logic [31:0] VFEQ_B             = 32'b1010000??????????011?????0110011;
  localparam logic [31:0] VFEQ_R_B           = 32'b1010000??????????111?????0110011;
  localparam logic [31:0] VFNE_B             = 32'b1010001??????????011?????0110011;
  localparam logic [31:0] VFNE_R_B           = 32'b1010001??????????111?????0110011;
  localparam logic [31:0] VFLT_B             = 32'b1010010??????????011?????0110011;
  localparam logic [31:0] VFLT_R_B           = 32'b1010010??????????111?????0110011;
  localparam logic [31:0] VFGE_B             = 32'b1010011??????????011?????0110011;
  localparam logic [31:0] VFGE_R_B           = 32'b1010011??????????111?????0110011;
  localparam logic [31:0] VFLE_B             = 32'b1010100??????????011?????0110011;
  localparam logic [31:0] VFLE_R_B           = 32'b1010100??????????111?????0110011;
  localparam logic [31:0] VFGT_B             = 32'b1010101??????????011?????0110011;
  localparam logic [31:0] VFGT_R_B           = 32'b1010101??????????111?????0110011;
  localparam logic [31:0] VFMV_X_B           = 32'b100110000000?????011?????0110011;
  localparam logic [31:0] VFMV_B_X           = 32'b100110000000?????111?????0110011;
  localparam logic [31:0] VFCLASS_B          = 32'b100110000001?????011?????0110011;
  localparam logic [31:0] VFCVT_X_B          = 32'b100110000010?????011?????0110011;
  localparam logic [31:0] VFCVT_XU_B         = 32'b100110000010?????111?????0110011;
  localparam logic [31:0] VFCVT_B_X          = 32'b100110000011?????011?????0110011;
  localparam logic [31:0] VFCVT_B_XU         = 32'b100110000011?????111?????0110011;
  localparam logic [31:0] VFCPKA_B_S         = 32'b1011000??????????011?????0110011;
  localparam logic [31:0] VFCPKB_B_S         = 32'b1011000??????????111?????0110011;
  localparam logic [31:0] VFCPKC_B_S         = 32'b1011001??????????011?????0110011;
  localparam logic [31:0] VFCPKD_B_S         = 32'b1011001??????????111?????0110011;
  localparam logic [31:0] VFCPKA_B_D         = 32'b1011010??????????011?????0110011;
  localparam logic [31:0] VFCPKB_B_D         = 32'b1011010??????????111?????0110011;
  localparam logic [31:0] VFCPKC_B_D         = 32'b1011011??????????011?????0110011;
  localparam logic [31:0] VFCPKD_B_D         = 32'b1011011??????????111?????0110011;
  localparam logic [31:0] VFCVT_S_B          = 32'b100110000111?????000?????0110011;
  localparam logic [31:0] VFCVTU_S_B         = 32'b100110000111?????100?????0110011;
  localparam logic [31:0] VFCVT_B_S          = 32'b100110000100?????011?????0110011;
  localparam logic [31:0] VFCVTU_B_S         = 32'b100110000100?????111?????0110011;
  localparam logic [31:0] VFCVT_H_B          = 32'b100110000111?????010?????0110011;
  localparam logic [31:0] VFCVTU_H_B         = 32'b100110000111?????110?????0110011;
  localparam logic [31:0] VFCVT_B_H          = 32'b100110000110?????011?????0110011;
  localparam logic [31:0] VFCVTU_B_H         = 32'b100110000110?????111?????0110011;
  localparam logic [31:0] VFCVT_AH_B         = 32'b100110000111?????001?????0110011;
  localparam logic [31:0] VFCVTU_AH_B        = 32'b100110000111?????101?????0110011;
  localparam logic [31:0] VFCVT_B_AH         = 32'b100110000101?????011?????0110011;
  localparam logic [31:0] VFCVTU_B_AH        = 32'b100110000101?????111?????0110011;
  localparam logic [31:0] VFDOTP_S           = 32'b1001010??????????000?????0110011;
  localparam logic [31:0] VFDOTP_R_S         = 32'b1001010??????????100?????0110011;
  localparam logic [31:0] VFAVG_S            = 32'b1010110??????????000?????0110011;
  localparam logic [31:0] VFAVG_R_S          = 32'b1010110??????????100?????0110011;
  localparam logic [31:0] FMULEX_S_H         = 32'b0100110??????????????????1010011;
  localparam logic [31:0] FMACEX_S_H         = 32'b0101010??????????????????1010011;
  localparam logic [31:0] VFDOTP_H           = 32'b1001010??????????010?????0110011;
  localparam logic [31:0] VFDOTP_R_H         = 32'b1001010??????????110?????0110011;
  localparam logic [31:0] VFDOTPEX_S_H       = 32'b1001011??????????010?????0110011;
  localparam logic [31:0] VFDOTPEX_S_R_H     = 32'b1001011??????????110?????0110011;
  localparam logic [31:0] VFAVG_H            = 32'b1010110??????????010?????0110011;
  localparam logic [31:0] VFAVG_R_H          = 32'b1010110??????????110?????0110011;
  localparam logic [31:0] FMULEX_S_AH        = 32'b0100110??????????101?????1010011;
  localparam logic [31:0] FMACEX_S_AH        = 32'b0101010??????????101?????1010011;
  localparam logic [31:0] VFDOTP_AH          = 32'b1001010??????????001?????0110011;
  localparam logic [31:0] VFDOTP_R_AH        = 32'b1001010??????????101?????0110011;
  localparam logic [31:0] VFDOTPEX_S_AH      = 32'b1001011??????????001?????0110011;
  localparam logic [31:0] VFDOTPEX_S_R_AH    = 32'b1001011??????????101?????0110011;
  localparam logic [31:0] VFAVG_AH           = 32'b1010110??????????001?????0110011;
  localparam logic [31:0] VFAVG_R_AH         = 32'b1010110??????????101?????0110011;
  localparam logic [31:0] FMULEX_S_B         = 32'b0100111??????????????????1010011;
  localparam logic [31:0] FMACEX_S_B         = 32'b0101011??????????????????1010011;
  localparam logic [31:0] VFDOTP_B           = 32'b1001010??????????011?????0110011;
  localparam logic [31:0] VFDOTP_R_B         = 32'b1001010??????????111?????0110011;
  localparam logic [31:0] VFDOTPEX_S_B       = 32'b1001011??????????011?????0110011;
  localparam logic [31:0] VFDOTPEX_S_R_B     = 32'b1001011??????????111?????0110011;
  localparam logic [31:0] VFAVG_B            = 32'b1010110??????????011?????0110011;
  localparam logic [31:0] VFAVG_R_B          = 32'b1010110??????????111?????0110011;
endpackage : fpu_ss_instr_pkg